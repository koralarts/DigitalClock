entity DigitalClock is

end DigitalClock;

architecture Behaviour of DigitalClock is

begin
end Behaviour;